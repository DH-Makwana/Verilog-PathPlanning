module node(add, o0, o1, o2, o3);
	input [4:0]add;
	output reg [0:6]o0, o1, o2, o3;
	
	reg [0:6]m[0:25][0:3];
	
	initial begin
	m[0][0] = {2'd3, 5'd1};
	m[0][1] = {2'd3, 5'd30};
	m[0][2] = {2'd3, 5'd30};
	m[0][3] = {2'd3, 5'd30};

	m[1][0] = {2'd3, 5'd0};
	m[1][1] = {2'd3, 5'd2};
	m[1][2] = {2'd3, 5'd13};
	m[1][3] = {2'd3, 5'd30};

	m[2][0] = {2'd3, 5'd1};
	m[2][1] = {2'd1, 5'd3};
	m[2][2] = {2'd3, 5'd5};
	m[2][3] = {2'd3, 5'd30};

	m[3][0] = {2'd1, 5'd2};
	m[3][1] = {2'd3, 5'd30};
	m[3][2] = {2'd3, 5'd30};
	m[3][3] = {2'd3, 5'd30};

	m[4][0] = {2'd3, 5'd6};
	m[4][1] = {2'd3, 5'd30};
	m[4][2] = {2'd3, 5'd30};
	m[4][3] = {2'd3, 5'd30};

	m[5][0] = {2'd3, 5'd2};
	m[5][1] = {2'd2, 5'd9};
	m[5][2] = {2'd1, 5'd6};
	m[5][3] = {2'd3, 5'd30};

	m[6][0] = {2'd3, 5'd4};
	m[6][1] = {2'd3, 5'd16};
	m[6][2] = {2'd1, 5'd5};
	m[6][3] = {2'd3, 5'd30};

	m[7][0] = {2'd2, 5'd12};
	m[7][1] = {2'd3, 5'd30};
	m[7][2] = {2'd3, 5'd30};
	m[7][3] = {2'd3, 5'd30};

	m[8][0] = {2'd1, 5'd9};
	m[8][1] = {2'd3, 5'd30};
	m[8][2] = {2'd3, 5'd30};
	m[8][3] = {2'd3, 5'd30};

	m[9][0] = {2'd1, 5'd8};
	m[9][1] = {2'd1, 5'd15};
	m[9][2] = {2'd2, 5'd5};
	m[9][3] = {2'd3, 5'd30};

	m[10][0] = {2'd2, 5'd16};
	m[10][1] = {2'd3, 5'd30};
	m[10][2] = {2'd3, 5'd30};
	m[10][3] = {2'd3, 5'd30};

	m[11][0] = {2'd3, 5'd12};
	m[11][1] = {2'd3, 5'd30};
	m[11][2] = {2'd3, 5'd30};
	m[11][3] = {2'd3, 5'd30};

	m[12][0] = {2'd3, 5'd11};
	m[12][1] = {2'd2, 5'd7};
	m[12][2] = {2'd1, 5'd13};
	m[12][3] = {2'd3, 5'd17};

	m[13][0] = {2'd1, 5'd12};
	m[13][1] = {2'd2, 5'd18};
	m[13][2] = {2'd3, 5'd1};
	m[13][3] = {2'd3, 5'd30};

	m[14][0] = {2'd1, 5'd15};
	m[14][1] = {2'd3, 5'd30};
	m[14][2] = {2'd3, 5'd30};
	m[14][3] = {2'd3, 5'd30};

	m[15][0] = {2'd1, 5'd14};
	m[15][1] = {2'd1, 5'd9};
	m[15][2] = {2'd1, 5'd22};
	m[15][3] = {2'd3, 5'd30};

	m[16][0] = {2'd2, 5'd10};
	m[16][1] = {2'd2, 5'd23};
	m[16][2] = {2'd3, 5'd6};
	m[16][3] = {2'd3, 5'd30};

	m[17][0] = {2'd3, 5'd12};
	m[17][1] = {2'd3, 5'd30};
	m[17][2] = {2'd3, 5'd30};
	m[17][3] = {2'd3, 5'd30};

	m[18][0] = {2'd1, 5'd19};
	m[18][1] = {2'd1, 5'd20};
	m[18][2] = {2'd2, 5'd13};
	m[18][3] = {2'd3, 5'd30};

	m[19][0] = {2'd1, 5'd18};
	m[19][1] = {2'd3, 5'd30};
	m[19][2] = {2'd3, 5'd30};
	m[19][3] = {2'd3, 5'd30};

	m[20][0] = {2'd1, 5'd18};
	m[20][1] = {2'd1, 5'd21};
	m[20][2] = {2'd2, 5'd22};
	m[20][3] = {2'd3, 5'd30};

	m[21][0] = {2'd1, 5'd20};
	m[21][1] = {2'd3, 5'd30};
	m[21][2] = {2'd3, 5'd30};
	m[21][3] = {2'd3, 5'd30};

	m[22][0] = {2'd1, 5'd23};
	m[22][1] = {2'd1, 5'd15};
	m[22][2] = {2'd2, 5'd20};
	m[22][3] = {2'd3, 5'd25};

	m[23][0] = {2'd1, 5'd22};
	m[23][1] = {2'd2, 5'd24};
	m[23][2] = {2'd2, 5'd16};
	m[23][3] = {2'd3, 5'd30};

	m[24][0] = {2'd2, 5'd23};
	m[24][1] = {2'd3, 5'd30};
	m[24][2] = {2'd3, 5'd30};
	m[24][3] = {2'd3, 5'd30};

	m[25][0] = {2'd3, 5'd22};
	m[25][1] = {2'd3, 5'd30};
	m[25][2] = {2'd3, 5'd30};
	m[25][3] = {2'd3, 5'd30};
	
	end
	always @(add)begin
		o0 = m[add][0];
		o1 = m[add][1];
		o2 = m[add][2];
		o3 = m[add][3];
	end
endmodule
